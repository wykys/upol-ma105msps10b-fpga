-------------------------------------------------------------------------------
-- ADC driver for AD9214
-- wykys 2020
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity adc_driver is
    generic (
        ADC_DATA_NUMBER_OF_BITS : positive := 10
    );
    port (
        -----------------------------------------------------------------------
        -- Clock --------------------------------------------------------------
        -----------------------------------------------------------------------
        clk_i : in std_logic;
        -----------------------------------------------------------------------
        -- Reset --------------------------------------------------------------
        -----------------------------------------------------------------------
        rst_i : in std_logic;
        -----------------------------------------------------------------------
        -- ADC interface ------------------------------------------------------
        -----------------------------------------------------------------------
        adc_ovrng_i : in std_logic;
        adc_data_i  : in std_logic_vector(ADC_DATA_NUMBER_OF_BITS - 1 downto 0);
        -----------------------------------------------------------------------
        -- Driver interface ---------------------------------------------------
        -----------------------------------------------------------------------
        adc_ovrng_o : out std_logic;
        adc_data_o  : out std_logic_vector(ADC_DATA_NUMBER_OF_BITS - 1 downto 0)
    );
end entity adc_driver;

architecture rtl of adc_driver is
begin

    ---------------------------------------------------------------------------
    -- Získání dat z ADC.
    ---------------------------------------------------------------------------
    process (clk_i) begin
        if rising_edge(clk_i) then
            if rst_i = '1' then
                ---------------------------------------------------------------
                -- Reset obvodu.
                ---------------------------------------------------------------
                adc_data_o  <= (others => '0');
                adc_ovrng_o <= '0';
            else
                ---------------------------------------------------------------
                -- Čtení dat z ADC.
                ---------------------------------------------------------------
                adc_data_o  <= adc_data_i;
                adc_ovrng_o <= adc_ovrng_i;
            end if;
        end if;
    end process;

end architecture rtl;